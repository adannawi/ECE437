/*
	Section for write back portion of pipeline

*/

module write_back (
	write_back_if.wb wbif
);


endmodule
