`include "caches_if.vh"
`include "cpu_types_pkg.vh"

module icache (
	caches_if.icache icif
	);

  // icache ports
  //dport icache (
  //  input   imemREN, imemaddr,
  //  output  ihit, imemload
  //);
  
endmodule