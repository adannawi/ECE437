
`include "cpu_types_pkg.vh"
`include "cache_control_if.vh"

module icache (
	caches_if.dcache icif
	);

endmodule