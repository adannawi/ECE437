`include "cache_control_if.vh"
`include "cpu_types_pkg.vh"

module icache (
	caches_if.icache icif
	);

endmodule