`include "hazard_unit_if.vh"
import cpu_types_pkg::*;

module hazard_unit
(
  input CLK, nRST,
  hazard_unit_if.hu huif
);
always_comb:
begin

end
endmodule
